module highScore ();









endmodule
